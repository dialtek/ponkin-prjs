// Create Date:    21:21:06 02/08/2014 
// Module Name:    m_seq_8bit 
//////////////////////////////////////////////////////////////////////////////////

module m_seq_8bit(						// ���������� ������ - �������� m_seq_8bit
  input clk,								// ������� �������� ������, ������� ������ � ����������
  output reg [7:0] LFSR = 1			// 8-������ ��������� �������, �������� �� ����. = 1
);

wire feedback = LFSR[7];				// "������" �������� �����, ������������ � �������� (8)
												// ���� ���������� �������� ���������� ����, 
												// �� ����� ����� �������� 8-�� ���� ���������� �������� - ��� �������� ������

always @(posedge clk)               // ��������� ���������������� �������� �� ��������� �������, ���-
                                    // ��������� �� ��������������(�����������) ������ ��������� �������

begin											// ������ ������

  LFSR[0] <= feedback;					// ������������ �������� ���� ���������� �������� �������� ����� 
												// �������� ����� (��������� �������� � �������� ����� ���������� ��������) 
  
  LFSR[1] <= LFSR[0];					// ������������ �������� 1-�� ���� -> 2-�� ����, ��� ����� 0-�� ���� � ������� �������
												// �������� �� 1 ���
												
  LFSR[2] <= LFSR[1];					// ������������ �������� 2-�� ���� -> 3-�� ����, ��� ����� 1-�� ���� � ������� �������
												// �������� �� 1 ���
  
  LFSR[3] <= LFSR[2];               // ������������ �������� 3-�� ���� -> 4-�� ����, ��� ����� 3-�� ���� � ������� �������
												// �������� �� 1 ���
  
  LFSR[4] <= LFSR[3] ^ feedback;    // ������������ 5-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 4-�� ����� �����. �������� � �������� �������� ����� (8-�� ��� �����. ��������)
											
  LFSR[5] <= LFSR[4] ^ feedback;    // ������������ 6-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 5-�� ����� �����. �������� � �������� �������� ����� (8-�� ��� �����. ��������)
  
  LFSR[6] <= LFSR[5] ^ feedback;    // ������������ 7-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 6-�� ����� �����. �������� � �������� �������� ����� (8-�� ��� �����. ��������)
  
  LFSR[7] <= LFSR[6];					// ������������ �������� 7-�� ���� -> 8-�� ����, ��� ����� 7-�� ���� � ������� �������
												// �������� �� 1 ���
												
end											// ����� ���������
endmodule	                        // ����� ��������� ������								


