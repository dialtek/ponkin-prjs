// Create Date:    21:21:06 02/08/2014 
// Module Name:    m_seq_8bit 
//////////////////////////////////////////////////////////////////////////////////

module m_seq_32bit(						// ���������� ������ - �������� m_seq_32bit
  input clk,								// ������� �������� ������, ������� ������ � ����������
  output reg [31:0] LFSR = 1			// 32-������ ��������� �������, �������� �� ����. = 1
);

wire feedback = LFSR[31];				// "������" �������� �����, ������������ � �������� (32)
												// ���� ���������� �������� ���������� ����, 
												// �� ����� ����� �������� 32-�� ���� ���������� �������� - ��� �������� ������

always @(posedge clk)               // ��������� ���������������� �������� �� ��������� �������, ���-
                                    // ��������� �� ��������������(�����������) ������ ��������� �������

begin											// ������ ������

  LFSR[0] <= feedback;					// ������������ �������� ���� ���������� �������� �������� ����� 
												// �������� ����� (��������� �������� � �������� ����� ���������� ��������) 
  
  LFSR[1]  <= LFSR[0];					// ����������� ����� ����� �������� �������� � ������� ������� ��������												
  LFSR[2]  <= LFSR[1];					
  LFSR[3]  <= LFSR[2];               
  LFSR[4]  <= LFSR[3];
  LFSR[5]  <= LFSR[4];															
  LFSR[6]  <= LFSR[5];					
  LFSR[7]  <= LFSR[6];               
  LFSR[8]  <= LFSR[7];
  LFSR[9]  <= LFSR[8];															
  LFSR[10] <= LFSR[9];					
  LFSR[11] <= LFSR[10];               
  LFSR[12] <= LFSR[11];
  LFSR[13] <= LFSR[12];															
  LFSR[14] <= LFSR[13];					
  LFSR[15] <= LFSR[14];               
  LFSR[16] <= LFSR[15];
  LFSR[17] <= LFSR[16];
  LFSR[18] <= LFSR[17];															
  LFSR[19] <= LFSR[18];					
  LFSR[20] <= LFSR[19];               
  LFSR[21] <= LFSR[20];
  LFSR[22] <= LFSR[21];															
  LFSR[23] <= LFSR[22];					
  LFSR[24] <= LFSR[23] ^ feedback;  // ������������ 25-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 24-�� ����� �����. �������� � �������� �������� ����� (32-�� ��� �����. ��������)		
  LFSR[25] <= LFSR[24] ^ feedback;	// ������������ 26-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 25-�� ����� �����. �������� � �������� �������� ����� (32-�� ��� �����. ��������)
  LFSR[26] <= LFSR[25];  
  LFSR[27] <= LFSR[26];					
  LFSR[28] <= LFSR[27];               
  LFSR[29] <= LFSR[28] ^ feedback;  // ������������ 30-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 29-�� ����� �����. �������� � �������� �������� ����� (32-�� ��� �����. ��������)
  LFSR[30] <= LFSR[29];															
  LFSR[31] <= LFSR[30] ^ feedback;	// ������������ 32-�� ���� �����. �������� ���������� �������� "������������ ��� (XOR)" 
											   // (�������� �� ������ "2") ����� 31-�� ����� �����. �������� � �������� �������� ����� (32-�� ��� �����. ��������)			            

end											// ����� ���������
endmodule	                        // ����� ��������� ������								


